// `define CFU_VERSION_13
// `define CFU_VERSION_12
// `define CFU_VERSION_11
`define CFU_VERSION_9
// `define CFU_VERSION_8
// `define CFU_VERSION_7
// `define CFU_VERSION_6
// `define CFU_VERSION_5
// `define CFU_VERSION_QUANT