// `define CFU_VERSION_14_1
// `define CFU_VERSION_14
// `define CFU_VERSION_13_2
// `define CFU_VERSION_13
// `define CFU_VERSION_12_3
// `define CFU_VERSION_12_2
// `define CFU_VERSION_12_1
`define CFU_VERSION_12_05
// `define CFU_VERSION_12
// `define CFU_VERSION_11_2
// `define CFU_VERSION_11_1
// `define CFU_VERSION_11
// `define CFU_VERSION_9
// `define CFU_VERSION_8
// `define CFU_VERSION_7
// `define CFU_VERSION_6
// `define CFU_VERSION_5
// `define CFU_VERSION_QUANT
// `define CFU_VERSION_9_TEST