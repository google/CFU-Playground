// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Rounding doubling high 32 bits. Given a 64 bit integer as {top, bottom}
// double and round to the nearest 2^32, outputting only the top half.

module rdh (
  // 64 bit integer as {top, bottom}
  input logic [31:0] top,
  input logic [31:0] bottom,

  output logic [31:0] out
);
  assign out = (signed'({top, bottom}) + 32'sh40000000) >> 31;
endmodule
